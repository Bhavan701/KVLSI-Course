// Code your design here
module jk_ff(j,k,clk,rst,q);
  input clk,rst,j,k;
  output q;
  reg temp;
  assign q=temp;
  always @ (posedge clk or posedge rst)
    begin
      if (rst)
        temp<=0;
      else 
        begin 
          if (j==0 && k==0)
            temp<=temp;
          else if (j==0 && k==0)
            temp<=0;
          else if (j==1 && k==0)
            temp<=1;
          else if (j==1&&k==1)
            temp<=~temp;
          else 
            temp<=temp;
        end 
    end
endmodule 