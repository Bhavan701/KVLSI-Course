// Code your design here
module xor_gate_w(output y, input a, input b);
  xor_gate my_xor(y, a, b);
endmodule