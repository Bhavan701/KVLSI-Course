// Code your design here

module xnor_gate_w(output y, input a, input b);
  xnor_gate my_xnor(y, a, b);
endmodule