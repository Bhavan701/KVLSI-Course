// Code your design here
// File: and_gate_udp.v
module and_gate_w(output y, input a, input b);
  and_gate my_and(y, a, b);
endmodule
