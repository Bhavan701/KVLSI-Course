// Code your design here
module or_gate_w(output y, input a, input b);
  or_gate my_or(y, a, b);
endmodule