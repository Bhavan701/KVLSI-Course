// Code your design here
module nand_gate_w(output y, input a, input b);
  nand_gate my_nand(y, a, b);
endmodule