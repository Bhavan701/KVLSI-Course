// Code your design here
 module nor_gate_w(output y, input a, input b);
  nor_gate my_nor(y, a, b);
endmodule