// Code your design here
module not_gate_w(output y, input a);
  not_gate my_not(y, a);
endmodule